`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/10/20 11:50:23
// Design Name: 
// Module Name: Shift
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Shift(A,Shift,EXT,Y,Z);
input [31:0] A;
input [4:0] Shift;
input EXT;
output [31:0] Y,Z;

reg [31:0] B,C,D;//SLL,SRL,SRA

always@(*) begin
case(Shift)
    5'b00000:B <= A;
    5'b00001:B <= {A[30:0],1'b0};
    5'b00010:B <= {A[29:0],2'b0};
    5'b00011:B <= {A[28:0],3'b0};
    5'b00100:B <= {A[27:0],4'b0};
    5'b00101:B <= {A[26:0],5'b0};
    5'b00110:B <= {A[25:0],6'b0};
    5'b00111:B <= {A[24:0],7'b0};
    5'b01000:B <= {A[23:0],8'b0};
    5'b01001:B <= {A[22:0],9'b0};
    5'b01010:B <= {A[21:0],10'b0};
    5'b01011:B <= {A[20:0],11'b0};
    5'b01100:B <= {A[19:0],12'b0};
    5'b01101:B <= {A[18:0],13'b0};
    5'b01110:B <= {A[17:0],14'b0};
    5'b01111:B <= {A[16:0],15'b0};
    5'b10000:B <= {A[15:0],16'b0};
    5'b10001:B <= {A[14:0],17'b0};
    5'b10010:B <= {A[13:0],18'b0};
    5'b10011:B <= {A[12:0],19'b0};
    5'b10100:B <= {A[11:0],20'b0};
    5'b10101:B <= {A[10:0],21'b0};
    5'b10110:B <= {A[9:0],22'b0};
    5'b10111:B <= {A[8:0],23'b0};
    5'b11000:B <= {A[7:0],24'b0};
    5'b11001:B <= {A[6:0],25'b0};
    5'b11010:B <= {A[5:0],26'b0};
    5'b11011:B <= {A[4:0],27'b0};
    5'b11100:B <= {A[3:0],28'b0};
    5'b11101:B <= {A[2:0],29'b0};
    5'b11110:B <= {A[1:0],30'b0};
    default:B <= {A[0],31'b0};
endcase

case(Shift)
    5'b00000:C <= A;
    5'b00001:C <= {1'b0,A[31:1]};
    5'b00010:C <= {2'b0,A[31:2]};
    5'b00011:C <= {3'b0,A[31:3]};
    5'b00100:C <= {4'b0,A[31:4]};
    5'b00101:C <= {5'b0,A[31:5]};
    5'b00110:C <= {6'b0,A[31:6]};
    5'b00111:C <= {7'b0,A[31:7]};
    5'b01000:C <= {8'b0,A[31:8]};
    5'b01001:C <= {9'b0,A[31:9]};
    5'b01010:C <= {10'b0,A[31:10]};
    5'b01011:C <= {11'b0,A[31:11]};
    5'b01100:C <= {12'b0,A[31:12]};
    5'b01101:C <= {13'b0,A[31:13]};
    5'b01110:C <= {14'b0,A[31:14]};
    5'b01111:C <= {15'b0,A[31:15]};
    5'b10000:C <= {16'b0,A[31:16]};
    5'b10001:C <= {17'b0,A[31:17]};
    5'b10010:C <= {18'b0,A[31:18]};
    5'b10011:C <= {19'b0,A[31:19]};
    5'b10100:C <= {20'b0,A[31:20]};
    5'b10101:C <= {21'b0,A[31:21]};
    5'b10110:C <= {22'b0,A[31:22]};
    5'b10111:C <= {23'b0,A[31:23]};
    5'b11000:C <= {24'b0,A[31:24]};
    5'b11001:C <= {25'b0,A[31:25]};
    5'b11010:C <= {26'b0,A[31:26]};
    5'b11011:C <= {27'b0,A[31:27]};
    5'b11100:C <= {28'b0,A[31:28]};
    5'b11101:C <= {29'b0,A[31:29]};
    5'b11110:C <= {30'b0,A[31:30]};
    default:C <= {31'b0,A[31]};
endcase

case(Shift)
    5'b00000:D <= A;
    5'b00001:D <= {1'h1,A[31:1]};
    5'b00010:D <= {2'h3,A[31:2]};
    5'b00011:D <= {3'h7,A[31:3]};
    5'b00100:D <= {4'hF,A[31:4]};
    5'b00101:D <= {5'h1F,A[31:5]};
    5'b00110:D <= {6'h3F,A[31:6]};
    5'b00111:D <= {7'h7F,A[31:7]};
    5'b01000:D <= {8'hFF,A[31:8]};
    5'b01001:D <= {9'h1FF,A[31:9]};
    5'b01010:D <= {10'h3FF,A[31:10]};
    5'b01011:D <= {11'h7FF,A[31:11]};
    5'b01100:D <= {12'hFFF,A[31:12]};
    5'b01101:D <= {13'h1FFF,A[31:13]};
    5'b01110:D <= {14'h3FFF,A[31:14]};
    5'b01111:D <= {15'h7FFF,A[31:15]};
    5'b10000:D <= {16'hFFFF,A[31:16]};
    5'b10001:D <= {17'h1FFFF,A[31:17]};
    5'b10010:D <= {18'h3FFFF,A[31:18]};
    5'b10011:D <= {19'h7FFFF,A[31:19]};
    5'b10100:D <= {20'hFFFFF,A[31:20]};
    5'b10101:D <= {21'h1FFFFF,A[31:21]};
    5'b10110:D <= {22'h3FFFFF,A[31:22]};
    5'b10111:D <= {23'h7FFFFF,A[31:23]};
    5'b11000:D <= {24'hFFFFFF,A[31:24]};
    5'b11001:D <= {25'h1FFFFFF,A[31:25]};
    5'b11010:D <= {26'h3FFFFFF,A[31:26]};
    5'b11011:D <= {27'h7FFFFFF,A[31:27]};
    5'b11100:D <= {28'hFFFFFFF,A[31:28]};
    5'b11101:D <= {29'h1FFFFFFF,A[31:29]};
    5'b11110:D <= {30'h3FFFFFFF,A[31:30]};
    default:D <= {31'h7FFFFFFF,A[31]};
endcase
end

assign Y = (EXT)?(A[31])?D:C:C;
assign Z = B;

endmodule
